package ahb_uvm_pkg;
 import uvm_pkg::*;
`include "uvm_macros.svh"
`include "amba_ahb_defines.v"
 `include "ahb_uvm_intf.sv"
 `include "ahb_uvm_seqitem.sv"
 `include "ahb_uvm_seq.sv"
 `include "ahb_uvm_sequencer.sv"
 `include "ahb_uvm_driver.sv"
 `include "ahb_uvm_monitor.sv"
 `include "ahb_uvm_agent.sv"
 `include "ahb_uvm_scoreboard.sv"
 `include "ahb_uvm_subscriber.sv"
 `include "ahb_uvm_env.sv"
 `include "ahb_uvm_test.sv"
endpackage: ahb_uvm_pkg